magic
tech scmos
timestamp 1749475690
<< nwell >>
rect 2 3 49 21
<< polysilicon >>
rect 9 13 11 15
rect 19 13 21 15
rect 29 13 31 15
rect 39 13 41 15
rect 9 -1 11 5
rect 19 -1 21 5
rect 29 -1 31 5
rect 9 -5 10 -1
rect 19 -5 20 -1
rect 29 -5 30 -1
rect 9 -16 11 -5
rect 19 -16 21 -5
rect 29 -16 31 -5
rect 39 -8 41 5
rect 40 -12 41 -8
rect 39 -16 41 -12
rect 9 -22 11 -20
rect 19 -22 21 -20
rect 29 -22 31 -20
rect 39 -22 41 -20
<< ndiffusion >>
rect 7 -20 9 -16
rect 11 -20 13 -16
rect 17 -20 19 -16
rect 21 -20 23 -16
rect 27 -20 29 -16
rect 31 -20 33 -16
rect 37 -20 39 -16
rect 41 -20 43 -16
<< pdiffusion >>
rect 3 9 9 13
rect 7 5 9 9
rect 11 5 19 13
rect 21 5 29 13
rect 31 9 33 13
rect 37 9 39 13
rect 31 5 39 9
rect 41 9 47 13
rect 41 5 43 9
<< metal1 >>
rect 6 17 10 21
rect 14 17 19 21
rect 23 17 27 21
rect 31 17 35 21
rect 39 17 44 21
rect 48 17 49 21
rect 33 13 37 17
rect 3 -8 7 5
rect 14 -5 16 -1
rect 24 -5 26 -1
rect 34 -5 36 -1
rect 43 -4 47 5
rect 43 -8 51 -4
rect 3 -12 36 -8
rect 3 -16 7 -12
rect 23 -16 27 -12
rect 43 -16 47 -8
rect 13 -24 17 -20
rect 33 -24 37 -20
rect 6 -28 10 -24
rect 14 -28 19 -24
rect 23 -28 27 -24
rect 31 -28 35 -24
rect 39 -28 44 -24
rect 48 -28 49 -24
<< ntransistor >>
rect 9 -20 11 -16
rect 19 -20 21 -16
rect 29 -20 31 -16
rect 39 -20 41 -16
<< ptransistor >>
rect 9 5 11 13
rect 19 5 21 13
rect 29 5 31 13
rect 39 5 41 13
<< polycontact >>
rect 10 -5 14 -1
rect 20 -5 24 -1
rect 30 -5 34 -1
rect 36 -12 40 -8
<< ndcontact >>
rect 3 -20 7 -16
rect 13 -20 17 -16
rect 23 -20 27 -16
rect 33 -20 37 -16
rect 43 -20 47 -16
<< pdcontact >>
rect 3 5 7 9
rect 33 9 37 13
rect 43 5 47 9
<< psubstratepcontact >>
rect 2 -28 6 -24
rect 10 -28 14 -24
rect 19 -28 23 -24
rect 27 -28 31 -24
rect 35 -28 39 -24
rect 44 -28 48 -24
<< nsubstratencontact >>
rect 2 17 6 21
rect 10 17 14 21
rect 19 17 23 21
rect 27 17 31 21
rect 35 17 39 21
rect 44 17 48 21
<< labels >>
rlabel metal1 36 -5 36 -1 7 in1
rlabel metal1 26 -5 26 -1 1 in2
rlabel metal1 16 -5 16 -1 1 in3
rlabel metal1 51 -8 51 -4 7 out
rlabel metal1 25 -26 25 -26 1 gnd!
rlabel metal1 25 19 25 19 5 vdd!
<< end >>
