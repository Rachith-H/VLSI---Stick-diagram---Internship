magic
tech scmos
timestamp 1749466325
<< nwell >>
rect 0 3 37 21
<< polysilicon >>
rect 8 13 10 15
rect 18 13 20 15
rect 28 13 30 15
rect 8 -1 10 5
rect 18 -1 20 5
rect 28 -1 30 5
rect 9 -5 10 -1
rect 19 -5 20 -1
rect 29 -5 30 -1
rect 8 -16 10 -5
rect 18 -16 20 -5
rect 28 -16 30 -5
rect 8 -22 10 -20
rect 18 -22 20 -20
rect 28 -22 30 -20
<< ndiffusion >>
rect 6 -20 8 -16
rect 10 -20 12 -16
rect 16 -20 18 -16
rect 20 -20 22 -16
rect 26 -20 28 -16
rect 30 -20 32 -16
<< pdiffusion >>
rect 6 9 8 13
rect 2 5 8 9
rect 10 5 18 13
rect 20 5 28 13
rect 30 9 36 13
rect 30 5 32 9
<< metal1 >>
rect 4 17 8 21
rect 12 17 16 21
rect 20 17 25 21
rect 29 17 33 21
rect 2 13 6 17
rect 3 -5 5 -1
rect 13 -5 15 -1
rect 23 -5 25 -1
rect 32 -8 36 5
rect 12 -12 39 -8
rect 12 -16 16 -12
rect 32 -16 36 -12
rect 2 -24 6 -20
rect 22 -24 26 -20
rect 4 -28 8 -24
rect 12 -28 16 -24
rect 20 -28 25 -24
rect 29 -28 33 -24
<< ntransistor >>
rect 8 -20 10 -16
rect 18 -20 20 -16
rect 28 -20 30 -16
<< ptransistor >>
rect 8 5 10 13
rect 18 5 20 13
rect 28 5 30 13
<< polycontact >>
rect 5 -5 9 -1
rect 15 -5 19 -1
rect 25 -5 29 -1
<< ndcontact >>
rect 2 -20 6 -16
rect 12 -20 16 -16
rect 22 -20 26 -16
rect 32 -20 36 -16
<< pdcontact >>
rect 2 9 6 13
rect 32 5 36 9
<< psubstratepcontact >>
rect 0 -28 4 -24
rect 8 -28 12 -24
rect 16 -28 20 -24
rect 25 -28 29 -24
rect 33 -28 37 -24
<< nsubstratencontact >>
rect 0 17 4 21
rect 8 17 12 21
rect 16 17 20 21
rect 25 17 29 21
rect 33 17 37 21
<< labels >>
rlabel metal1 22 19 22 19 5 vdd!
rlabel metal1 22 -26 22 -26 1 gnd!
rlabel metal1 3 -5 3 -1 3 in1
rlabel metal1 13 -5 13 -1 1 in2
rlabel metal1 23 -5 23 -1 1 in3
rlabel metal1 39 -12 39 -8 7 out
<< end >>
