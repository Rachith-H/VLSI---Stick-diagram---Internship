magic
tech scmos
timestamp 1749467560
<< nwell >>
rect -3 1 47 19
<< polysilicon >>
rect 6 11 8 13
rect 16 11 18 13
rect 26 11 28 13
rect 36 11 38 13
rect 6 -16 8 3
rect 16 -16 18 3
rect 26 -16 28 3
rect 36 -7 38 3
rect 37 -11 38 -7
rect 6 -20 7 -16
rect 16 -20 17 -16
rect 26 -20 27 -16
rect 6 -25 8 -20
rect 16 -25 18 -20
rect 26 -25 28 -20
rect 36 -25 38 -11
rect 6 -31 8 -29
rect 16 -31 18 -29
rect 26 -31 28 -29
rect 36 -31 38 -29
<< ndiffusion >>
rect 3 -29 6 -25
rect 8 -29 16 -25
rect 18 -29 26 -25
rect 28 -29 30 -25
rect 34 -29 36 -25
rect 38 -29 41 -25
<< pdiffusion >>
rect -1 7 6 11
rect 3 3 6 7
rect 8 7 10 11
rect 14 7 16 11
rect 8 3 16 7
rect 18 7 26 11
rect 18 3 20 7
rect 24 3 26 7
rect 28 7 30 11
rect 34 7 36 11
rect 28 3 36 7
rect 38 7 45 11
rect 38 3 41 7
<< metal1 >>
rect 1 15 5 19
rect 9 15 15 19
rect 19 15 24 19
rect 28 15 32 19
rect 36 15 41 19
rect 10 11 14 15
rect 30 11 34 15
rect -1 -7 3 3
rect 20 -7 24 3
rect 41 -7 45 3
rect -1 -11 33 -7
rect 41 -11 48 -7
rect -1 -25 3 -11
rect 11 -20 14 -16
rect 21 -20 24 -16
rect 31 -20 34 -16
rect 41 -25 45 -11
rect 30 -33 34 -29
rect 1 -37 5 -33
rect 9 -37 15 -33
rect 19 -37 24 -33
rect 28 -37 32 -33
rect 36 -37 41 -33
<< ntransistor >>
rect 6 -29 8 -25
rect 16 -29 18 -25
rect 26 -29 28 -25
rect 36 -29 38 -25
<< ptransistor >>
rect 6 3 8 11
rect 16 3 18 11
rect 26 3 28 11
rect 36 3 38 11
<< polycontact >>
rect 33 -11 37 -7
rect 7 -20 11 -16
rect 17 -20 21 -16
rect 27 -20 31 -16
<< ndcontact >>
rect -1 -29 3 -25
rect 30 -29 34 -25
rect 41 -29 45 -25
<< pdcontact >>
rect -1 3 3 7
rect 10 7 14 11
rect 20 3 24 7
rect 30 7 34 11
rect 41 3 45 7
<< psubstratepcontact >>
rect -3 -37 1 -33
rect 5 -37 9 -33
rect 15 -37 19 -33
rect 24 -37 28 -33
rect 32 -37 36 -33
rect 41 -37 45 -33
<< nsubstratencontact >>
rect -3 15 1 19
rect 5 15 9 19
rect 15 15 19 19
rect 24 15 28 19
rect 32 15 36 19
rect 41 15 45 19
<< labels >>
rlabel metal1 14 -20 14 -16 1 in3
rlabel metal1 24 -20 24 -16 1 in2
rlabel metal1 34 -20 34 -16 7 in1
rlabel metal1 12 -35 12 -35 1 gnd!
rlabel metal1 12 17 12 17 5 vdd!
rlabel metal1 48 -11 48 -7 7 out
<< end >>
