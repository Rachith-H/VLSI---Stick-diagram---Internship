* SPICE3 file created from or2.ext - technology: scmos

.model pfet pmos (LEVEL=1 VTO=-0.7 KP=25u LAMBDA=0.02)
.model nfet nmos (LEVEL=1 VTO=0.7 KP=50u LAMBDA=0.02)

.option scale=1u

M1000 out a_22_5# gnd Gnd nfet w=4 l=2
+  ad=24p pd=20u as=16p ps=12u
M1001 gnd in1 a_22_5# Gnd nfet w=4 l=2
+  ad=16p pd=12u as=16p ps=12u
M1002 a_22_5# in2 a_22_5# Gnd nfet w=4 l=2
+  ad=28p pd=22u as=60p ps=46u
M1003 a_31_29# in2 a_22_5# vdd pfet w=8 l=2
+  ad=32p pd=16u as=56p ps=30u
M1004 vdd in1 a_31_29# vdd pfet w=8 l=2
+  ad=32p pd=16u as=32p ps=16u
M1005 out a_22_5# vdd vdd pfet w=8 l=2
+  ad=48p pd=28u as=32p ps=16u
C0 out 0 4.136f 
C1 a_22_5# 0 14.53f 
C2 in1 0 7.684f 
C3 in2 0 7.684f 

v1 vdd gnd 1.8
vina in1 gnd pulse(0 1.8 0n 1n 1n 50n 100n)
vinb in2 gnd pulse(0 1.8 0n 1n 1n 100n 200n)

.tran 1n 400n
.control
run 
plot v(in1)+2 v(in2)+4 v(out)
.endc
.end
