magic
tech scmos
timestamp 1749364935
<< nwell >>
rect -3 1 36 19
<< polysilicon >>
rect 5 11 7 13
rect 15 11 17 13
rect 25 11 27 13
rect 5 -16 7 3
rect 15 -16 17 3
rect 25 -16 27 3
rect 6 -20 7 -16
rect 16 -20 17 -16
rect 26 -20 27 -16
rect 5 -25 7 -20
rect 15 -25 17 -20
rect 25 -25 27 -20
rect 5 -31 7 -29
rect 15 -31 17 -29
rect 25 -31 27 -29
<< ndiffusion >>
rect 3 -29 5 -25
rect 7 -29 15 -25
rect 17 -29 25 -25
rect 27 -29 30 -25
<< pdiffusion >>
rect 3 7 5 11
rect -1 3 5 7
rect 7 7 15 11
rect 7 3 9 7
rect 13 3 15 7
rect 17 7 19 11
rect 23 7 25 11
rect 17 3 25 7
rect 27 7 34 11
rect 27 3 30 7
<< metal1 >>
rect 1 15 5 19
rect 9 15 14 19
rect 18 15 24 19
rect 28 15 32 19
rect -1 11 3 15
rect 19 11 23 15
rect 9 -7 13 3
rect 30 -7 34 3
rect 9 -11 37 -7
rect -1 -20 2 -16
rect 9 -20 12 -16
rect 19 -20 22 -16
rect 30 -25 34 -11
rect -1 -33 3 -29
rect 1 -37 5 -33
rect 9 -37 14 -33
rect 18 -37 24 -33
rect 28 -37 32 -33
<< ntransistor >>
rect 5 -29 7 -25
rect 15 -29 17 -25
rect 25 -29 27 -25
<< ptransistor >>
rect 5 3 7 11
rect 15 3 17 11
rect 25 3 27 11
<< polycontact >>
rect 2 -20 6 -16
rect 12 -20 16 -16
rect 22 -20 26 -16
<< ndcontact >>
rect -1 -29 3 -25
rect 30 -29 34 -25
<< pdcontact >>
rect -1 7 3 11
rect 9 3 13 7
rect 19 7 23 11
rect 30 3 34 7
<< psubstratepcontact >>
rect -3 -37 1 -33
rect 5 -37 9 -33
rect 14 -37 18 -33
rect 24 -37 28 -33
rect 32 -37 36 -33
<< nsubstratencontact >>
rect -3 15 1 19
rect 5 15 9 19
rect 14 15 18 19
rect 24 15 28 19
rect 32 15 36 19
<< labels >>
rlabel metal1 21 17 21 17 5 vdd!
rlabel metal1 21 -35 21 -35 1 gnd!
rlabel metal1 -1 -20 -1 -16 3 in1
rlabel metal1 9 -20 9 -16 1 in2
rlabel metal1 19 -20 19 -16 1 in3
rlabel metal1 37 -11 37 -7 7 out
<< end >>
