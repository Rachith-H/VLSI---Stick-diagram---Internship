* SPICE3 file created from nand2.ext - technology: scmos


.model pfet pmos (LEVEL=1 VTO=-0.7 KP=25u LAMBDA=0.02)
.model nfet nmos (LEVEL=1 VTO=0.7 KP=50u LAMBDA=0.02)


.option scale=1u

M1000 gnd in2 a_4_n28# Gnd nfet w=4 l=2
+  ad=24p pd=20u as=20p ps=14u
M1001 vdd in2 out vdd pfet w=8 l=2
+  ad=48p pd=28u as=40p ps=18u
M1002 a_4_n28# in1 out Gnd nfet w=4 l=2
+  ad=20p pd=14u as=24p ps=20u
M1003 out in1 vdd vdd pfet w=8 l=2
+  ad=40p pd=18u as=48p ps=28u
C0 out 0 8.272f 
C1 in2 0 9.498f 
C2 in1 0 9.626f 


v1 vdd gnd 1.8
vina in1 gnd pulse(0 1.8 0n 1n 1n 50n 100n)
vinb in2 gnd pulse(0 1.8 0n 1n 1n 100n 200n)

.tran 1n 400n
.control
run 
plot v(in1)+2 v(in2)+4 v(out)
.endc
.end
