magic
tech scmos
timestamp 1749131706
<< nwell >>
rect -9 26 13 48
<< polysilicon >>
rect 1 38 3 40
rect 1 19 3 30
rect 2 14 3 19
rect 1 4 3 14
rect 1 -2 3 0
<< ndiffusion >>
rect -1 0 1 4
rect 3 0 5 4
<< pdiffusion >>
rect -1 34 1 38
rect -5 30 1 34
rect 3 34 9 38
rect 3 30 5 34
<< metal1 >>
rect -4 43 0 47
rect 4 43 8 47
rect -8 42 12 43
rect -5 38 -1 42
rect 5 19 9 30
rect -11 14 -2 19
rect 5 15 16 19
rect 5 4 9 15
rect -5 -6 -1 0
rect -4 -10 0 -6
rect 4 -10 8 -6
<< ntransistor >>
rect 1 0 3 4
<< ptransistor >>
rect 1 30 3 38
<< polycontact >>
rect -2 14 2 19
<< ndcontact >>
rect -5 0 -1 4
rect 5 0 9 4
<< pdcontact >>
rect -5 34 -1 38
rect 5 30 9 34
<< psubstratepcontact >>
rect -8 -10 -4 -6
rect 0 -10 4 -6
rect 8 -10 12 -6
<< nsubstratencontact >>
rect -8 43 -4 47
rect 0 43 4 47
rect 8 43 12 47
<< labels >>
rlabel metal1 6 -8 6 -8 1 gnd!
rlabel metal1 -2 45 -2 45 5 vdd!
rlabel metal1 -11 14 -11 19 3 in
rlabel metal1 16 15 16 19 7 out
<< end >>
