magic
tech scmos
timestamp 1749706281
<< nwell >>
rect -9 26 61 47
<< polysilicon >>
rect 1 38 3 40
rect 25 38 27 40
rect 49 38 51 40
rect 1 19 3 30
rect 25 19 27 30
rect 49 19 51 30
rect 2 15 3 19
rect 26 15 27 19
rect 50 15 51 19
rect 1 4 3 15
rect 25 4 27 15
rect 49 4 51 15
rect 1 -2 3 0
rect 25 -2 27 0
rect 49 -2 51 0
<< ndiffusion >>
rect -1 0 1 4
rect 3 0 5 4
rect 23 0 25 4
rect 27 0 29 4
rect 47 0 49 4
rect 51 0 53 4
<< pdiffusion >>
rect -1 34 1 38
rect -5 30 1 34
rect 3 34 9 38
rect 3 30 5 34
rect 23 34 25 38
rect 19 30 25 34
rect 27 34 33 38
rect 27 30 29 34
rect 47 34 49 38
rect 43 30 49 34
rect 51 34 57 38
rect 51 30 53 34
<< metal1 >>
rect -4 43 0 47
rect 4 43 8 47
rect 12 43 16 47
rect 20 43 24 47
rect 28 43 32 47
rect 36 43 40 47
rect 44 43 48 47
rect 52 43 56 47
rect -5 38 -1 43
rect 19 38 23 43
rect 43 38 47 43
rect 5 19 9 30
rect 29 19 33 30
rect 53 19 57 30
rect -15 15 -2 19
rect 5 15 22 19
rect 29 15 46 19
rect 53 15 70 19
rect -15 -13 -11 15
rect 5 4 9 15
rect 29 4 33 15
rect 53 4 57 15
rect -5 -6 -1 0
rect 19 -6 23 0
rect 43 -6 47 0
rect -4 -10 0 -6
rect 4 -10 8 -6
rect 12 -10 16 -6
rect 20 -10 24 -6
rect 28 -10 32 -6
rect 36 -10 40 -6
rect 44 -10 48 -6
rect 52 -10 56 -6
rect 63 -13 67 15
rect -15 -17 67 -13
<< ntransistor >>
rect 1 0 3 4
rect 25 0 27 4
rect 49 0 51 4
<< ptransistor >>
rect 1 30 3 38
rect 25 30 27 38
rect 49 30 51 38
<< polycontact >>
rect -2 15 2 19
rect 22 15 26 19
rect 46 15 50 19
<< ndcontact >>
rect -5 0 -1 4
rect 5 0 9 4
rect 19 0 23 4
rect 29 0 33 4
rect 43 0 47 4
rect 53 0 57 4
<< pdcontact >>
rect -5 34 -1 38
rect 5 30 9 34
rect 19 34 23 38
rect 29 30 33 34
rect 43 34 47 38
rect 53 30 57 34
<< psubstratepcontact >>
rect -8 -10 -4 -6
rect 0 -10 4 -6
rect 8 -10 12 -6
rect 16 -10 20 -6
rect 24 -10 28 -6
rect 32 -10 36 -6
rect 40 -10 44 -6
rect 48 -10 52 -6
rect 56 -10 60 -6
<< nsubstratencontact >>
rect -8 43 -4 47
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
rect 32 43 36 47
rect 40 43 44 47
rect 48 43 52 47
rect 56 43 60 47
<< labels >>
rlabel metal1 30 45 30 45 5 vdd!
rlabel metal1 30 -8 30 -8 1 gnd!
rlabel metal1 70 15 70 19 7 out
<< end >>
