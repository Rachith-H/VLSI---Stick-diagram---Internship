magic
tech scmos
timestamp 1749293991
<< nwell >>
rect -4 6 28 25
<< polysilicon >>
rect 5 16 7 18
rect 17 16 19 18
rect 5 2 7 8
rect 17 2 19 8
rect 6 -2 7 2
rect 18 -2 19 2
rect 5 -18 7 -2
rect 17 -18 19 -2
rect 5 -24 7 -22
rect 17 -24 19 -22
<< ndiffusion >>
rect 2 -22 5 -18
rect 7 -22 10 -18
rect 14 -22 17 -18
rect 19 -22 22 -18
<< pdiffusion >>
rect 2 12 5 16
rect -2 8 5 12
rect 7 8 17 16
rect 19 12 26 16
rect 19 8 22 12
<< metal1 >>
rect 0 21 4 25
rect 8 21 16 25
rect 20 21 24 25
rect -2 16 2 21
rect -2 -2 2 2
rect 10 -2 14 2
rect 22 -8 26 8
rect -2 -12 30 -8
rect -2 -18 2 -12
rect 22 -18 26 -12
rect 10 -28 14 -22
rect 0 -32 4 -28
rect 8 -32 16 -28
rect 20 -32 24 -28
<< ntransistor >>
rect 5 -22 7 -18
rect 17 -22 19 -18
<< ptransistor >>
rect 5 8 7 16
rect 17 8 19 16
<< polycontact >>
rect 2 -2 6 2
rect 14 -2 18 2
<< ndcontact >>
rect -2 -22 2 -18
rect 10 -22 14 -18
rect 22 -22 26 -18
<< pdcontact >>
rect -2 12 2 16
rect 22 8 26 12
<< psubstratepcontact >>
rect -4 -32 0 -28
rect 4 -32 8 -28
rect 16 -32 20 -28
rect 24 -32 28 -28
<< nsubstratencontact >>
rect -4 21 0 25
rect 4 21 8 25
rect 16 21 20 25
rect 24 21 28 25
<< labels >>
rlabel metal1 12 -30 12 -30 1 gnd!
rlabel metal1 12 23 12 23 5 vdd!
rlabel metal1 -2 -2 -2 2 3 in1
rlabel metal1 10 -2 10 2 1 in2
rlabel metal1 30 -12 30 -8 7 out
<< end >>
