* SPICE3 file created from /home/rachith/Desktop/Layouts/nor2.ext - technology: scmos

.model pfet pmos (LEVEL=1 VTO=-0.7 KP=25u LAMBDA=0.02)
.model nfet nmos (LEVEL=1 VTO=0.7 KP=50u LAMBDA=0.02)

.option scale=1u

M1000 a_7_8# in1 vdd vdd pfet w=8 l=2
+  ad=40p pd=18u as=56p ps=30u
M1001 out in2 gnd Gnd nfet w=4 l=2
+  ad=28p pd=22u as=20p ps=14u
M1002 out in2 a_7_8# vdd pfet w=8 l=2
+  ad=56p pd=30u as=40p ps=18u
M1003 gnd in1 out Gnd nfet w=4 l=2
+  ad=20p pd=14u as=28p ps=22u
C0 out 0 10.152f 
C1 in2 0 9.488f 
C2 in1 0 9.488f 

v1 vdd gnd 1.8
vina in1 gnd pulse(0 1.8 0n 1n 1n 50n 100n)
vinb in2 gnd pulse(0 1.8 0n 1n 1n 100n 200n)

.tran 1n 400n
.control
run 
plot v(in1)+2 v(in2)+4 v(out)
.endc
.end
