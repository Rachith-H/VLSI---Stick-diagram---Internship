magic
tech scmos
timestamp 1749826122
<< nwell >>
rect -49 8 68 33
<< polysilicon >>
rect -39 18 -37 20
rect -29 18 -27 20
rect -19 18 -17 20
rect -1 18 1 20
rect 9 18 11 20
rect 27 18 29 20
rect 37 18 39 20
rect 47 18 49 20
rect 57 18 59 20
rect -39 -21 -37 10
rect -29 -7 -27 10
rect -28 -11 -27 -7
rect -39 -25 -38 -21
rect -39 -45 -37 -25
rect -29 -45 -27 -11
rect -19 -7 -17 10
rect -19 -11 -18 -7
rect -19 -45 -17 -11
rect -1 -15 1 10
rect 9 -7 11 10
rect 27 -7 29 10
rect 9 -11 10 -7
rect -1 -19 0 -15
rect -1 -45 1 -19
rect 9 -45 11 -11
rect 27 -45 29 -11
rect 37 -15 39 10
rect 37 -45 39 -19
rect 47 -22 49 10
rect 57 0 59 10
rect 58 -4 59 0
rect 48 -26 49 -22
rect 47 -45 49 -26
rect 57 -29 59 -4
rect 58 -33 59 -29
rect 57 -45 59 -33
rect -39 -52 -37 -49
rect -29 -51 -27 -49
rect -19 -51 -17 -49
rect -1 -51 1 -49
rect 9 -51 11 -49
rect 27 -51 29 -49
rect 37 -51 39 -49
rect 47 -51 49 -49
rect 57 -51 59 -49
<< ndiffusion >>
rect -41 -49 -39 -45
rect -37 -49 -35 -45
rect -31 -49 -29 -45
rect -27 -49 -19 -45
rect -17 -49 -15 -45
rect -3 -49 -1 -45
rect 1 -49 3 -45
rect 7 -49 9 -45
rect 11 -49 13 -45
rect 25 -49 27 -45
rect 29 -49 37 -45
rect 39 -49 41 -45
rect 45 -49 47 -45
rect 49 -49 57 -45
rect 59 -49 62 -45
<< pdiffusion >>
rect -45 14 -39 18
rect -41 10 -39 14
rect -37 14 -35 18
rect -31 14 -29 18
rect -37 10 -29 14
rect -27 14 -19 18
rect -27 10 -25 14
rect -21 10 -19 14
rect -17 14 -15 18
rect -17 10 -11 14
rect -7 14 -1 18
rect -3 10 -1 14
rect 1 14 3 18
rect 7 14 9 18
rect 1 10 9 14
rect 11 14 17 18
rect 11 10 13 14
rect 21 14 27 18
rect 25 10 27 14
rect 29 14 31 18
rect 35 14 37 18
rect 29 10 37 14
rect 39 14 47 18
rect 39 10 41 14
rect 45 10 47 14
rect 49 14 51 18
rect 55 14 57 18
rect 49 10 57 14
rect 59 14 66 18
rect 59 10 62 14
<< metal1 >>
rect -45 29 -41 33
rect -37 29 -33 33
rect -29 29 -25 33
rect -21 29 -17 33
rect -13 29 -9 33
rect -5 29 -1 33
rect -35 18 -31 29
rect -15 18 -11 29
rect 3 18 7 33
rect 11 29 15 33
rect 19 29 23 33
rect 27 29 32 33
rect 36 29 40 33
rect 44 29 48 33
rect 52 29 56 33
rect 60 29 64 33
rect 31 18 35 29
rect 51 22 74 26
rect 51 18 55 22
rect -45 -13 -41 10
rect -35 -11 -32 -7
rect -51 -17 -41 -13
rect -45 -45 -41 -17
rect -25 -21 -21 10
rect -14 -11 -11 -7
rect -34 -25 -11 -21
rect -15 -45 -11 -25
rect -7 -22 -3 10
rect 13 0 17 10
rect 21 7 25 10
rect 41 7 45 10
rect 62 7 66 10
rect 21 3 66 7
rect 13 -4 54 0
rect 14 -11 25 -7
rect 29 -11 31 -7
rect 70 -10 74 22
rect 66 -14 74 -10
rect 4 -19 35 -15
rect 39 -19 41 -15
rect -7 -26 44 -22
rect -7 -45 -3 -26
rect 13 -33 54 -29
rect 13 -45 17 -33
rect 70 -36 74 -14
rect 21 -40 74 -36
rect 21 -45 25 -40
rect 62 -45 66 -40
rect -35 -54 -31 -49
rect -45 -58 -41 -54
rect -37 -58 -33 -54
rect -29 -58 -25 -54
rect -21 -58 -17 -54
rect -13 -58 -9 -54
rect -5 -58 -1 -54
rect 3 -58 7 -49
rect 41 -54 45 -49
rect 11 -58 15 -54
rect 19 -58 24 -54
rect 28 -58 32 -54
rect 36 -58 40 -54
rect 44 -58 48 -54
rect 52 -58 56 -54
rect 60 -58 64 -54
<< ntransistor >>
rect -39 -49 -37 -45
rect -29 -49 -27 -45
rect -19 -49 -17 -45
rect -1 -49 1 -45
rect 9 -49 11 -45
rect 27 -49 29 -45
rect 37 -49 39 -45
rect 47 -49 49 -45
rect 57 -49 59 -45
<< ptransistor >>
rect -39 10 -37 18
rect -29 10 -27 18
rect -19 10 -17 18
rect -1 10 1 18
rect 9 10 11 18
rect 27 10 29 18
rect 37 10 39 18
rect 47 10 49 18
rect 57 10 59 18
<< polycontact >>
rect -32 -11 -28 -7
rect -38 -25 -34 -21
rect -18 -11 -14 -7
rect 10 -11 14 -7
rect 25 -11 29 -7
rect 0 -19 4 -15
rect 35 -19 39 -15
rect 54 -4 58 0
rect 44 -26 48 -22
rect 54 -33 58 -29
<< ndcontact >>
rect -45 -49 -41 -45
rect -35 -49 -31 -45
rect -15 -49 -11 -45
rect -7 -49 -3 -45
rect 3 -49 7 -45
rect 13 -49 17 -45
rect 21 -49 25 -45
rect 41 -49 45 -45
rect 62 -49 66 -45
<< pdcontact >>
rect -45 10 -41 14
rect -35 14 -31 18
rect -25 10 -21 14
rect -15 14 -11 18
rect -7 10 -3 14
rect 3 14 7 18
rect 13 10 17 14
rect 21 10 25 14
rect 31 14 35 18
rect 41 10 45 14
rect 51 14 55 18
rect 62 10 66 14
<< psubstratepcontact >>
rect -49 -58 -45 -54
rect -41 -58 -37 -54
rect -33 -58 -29 -54
rect -25 -58 -21 -54
rect -17 -58 -13 -54
rect -9 -58 -5 -54
rect -1 -58 3 -54
rect 7 -58 11 -54
rect 15 -58 19 -54
rect 24 -58 28 -54
rect 32 -58 36 -54
rect 40 -58 44 -54
rect 48 -58 52 -54
rect 56 -58 60 -54
rect 64 -58 68 -54
<< nsubstratencontact >>
rect -49 29 -45 33
rect -41 29 -37 33
rect -33 29 -29 33
rect -25 29 -21 33
rect -17 29 -13 33
rect -9 29 -5 33
rect -1 29 3 33
rect 7 29 11 33
rect 15 29 19 33
rect 23 29 27 33
rect 32 29 36 33
rect 40 29 44 33
rect 48 29 52 33
rect 56 29 60 33
rect 64 29 68 33
<< labels >>
rlabel metal1 31 -11 31 -7 1 in1
rlabel metal1 41 -19 41 -15 1 in2
rlabel metal1 30 -56 30 -56 1 gnd!
rlabel metal1 30 31 30 31 5 vdd!
rlabel metal1 -11 -11 -11 -7 1 in1
rlabel metal1 -35 -11 -35 -7 1 in2
rlabel metal1 66 -14 66 -10 1 sum
rlabel metal1 -51 -17 -51 -13 3 carry
<< end >>
